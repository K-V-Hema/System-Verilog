module tb;
int arr[][][];
int i,j,k;
initial begin
		arr=new[5];
	for(i=0;i<5;i++)begin
		arr[i]=new[4];
	for(j=0;j<4;j++)begin
		arr[i][j]=new[3];
	for(k=0;k<2;k++)begin
		arr[i][j][k]=$urandom_range(10,100);
	end
	end
	end
$display("arr=%p",arr);
end
endmodule

/*arr='{'{'{73, 67, 67}, '{83, 86, 27}, '{38, 80, 47}, '{51, 59, 43}},
		'{'{65, 43, 53}, '{57, 39, 66}, '{25, 71, 64}, '{17, 43, 79}},
		'{'{55, 44, 59}, '{95, 33, 94}, '{35, 71, 82}, '{83, 24, 82}},
		'{'{27, 91, 14}, '{39, 89, 45}, '{74, 71, 95}, '{68, 10, 19}},
		'{'{75, 14, 58}, '{71, 38, 92}, '{91, 73, 63}, '{34, 59, 60}}}*/
